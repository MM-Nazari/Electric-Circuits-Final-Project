** Profile: "SCHEMATIC1-FinalProject-Part2"  [ x:\orcad\capture\finalproject-mmnazari-9931061\finalproject-part2\simulation\finalproject-part2-schematic1-finalproject-part2.sim ] 

** Creating circuit file "finalproject-part2-schematic1-finalproject-part2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10k 0.001 10k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\finalproject-part2-SCHEMATIC1.net" 


.END
