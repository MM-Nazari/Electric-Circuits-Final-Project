** Profile: "SCHEMATIC1-FinalProject-Part3"  [ x:\orcad\capture\finalproject-mmnazari-9931061\finalproject-part3\simulation\finalproject-part3-schematic1-finalproject-part3.sim ] 

** Creating circuit file "finalproject-part3-schematic1-finalproject-part3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10k 0.001 10k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\finalproject-part3-SCHEMATIC1.net" 


.END
