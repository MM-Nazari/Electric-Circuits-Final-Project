** Profile: "SCHEMATIC1-FinalProject-Part6-Vth"  [ x:\orcad\capture\finalproject-mmnazari-9931061\finalproject-part6\simulation\vth\finalproject-part6-vth-schematic1-finalproject-part6-vth.sim ] 

** Creating circuit file "finalproject-part6-vth-schematic1-finalproject-part6-vth.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1 0.318 0.318
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\finalproject-part6-vth-SCHEMATIC1.net" 


.END
