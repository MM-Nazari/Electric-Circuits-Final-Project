** Profile: "SCHEMATIC1-FinalProject-Part1"  [ x:\orcad\capture\finalproject-mmnazari-9931061\finalproject-part1\simulation\finalproject-part1-schematic1-finalproject-part1.sim ] 

** Creating circuit file "finalproject-part1-schematic1-finalproject-part1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 15.707 0 15.707m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\finalproject-part1-SCHEMATIC1.net" 


.END
