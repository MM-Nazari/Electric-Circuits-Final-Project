** Profile: "SCHEMATIC1-FinalProject-Part4"  [ x:\orcad\capture\finalproject-mmnazari-9931061\finalproject-part4\simulation\finalproject-part4-schematic1-finalproject-part4.sim ] 

** Creating circuit file "finalproject-part4-schematic1-finalproject-part4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM C9 10n 500n 1n 
+ LIN V_V17 0.01 -0.01 -0.001 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\finalproject-part4-SCHEMATIC1.net" 


.END
